
module test(
	input wire foo,
	output wire bar
);

	assign foo = bar;

endmodule
